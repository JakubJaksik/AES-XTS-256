module AesSboxFun (
	input	wire	[7:0]	inData,	
    output	wire	[7:0]	outData 
);


assign outData = 	(inData == 8'h00) ? 8'h63 :
					(inData == 8'h01) ? 8'h7C :
					(inData == 8'h02) ? 8'h77 :
					(inData == 8'h03) ? 8'h7B :
					(inData == 8'h04) ? 8'hF2 :
					(inData == 8'h05) ? 8'h6B :
					(inData == 8'h06) ? 8'h6F :
					(inData == 8'h07) ? 8'hC5 :
					(inData == 8'h08) ? 8'h30 :
					(inData == 8'h09) ? 8'h01 :
					(inData == 8'h0A) ? 8'h67 :
					(inData == 8'h0B) ? 8'h2B :
					(inData == 8'h0C) ? 8'hFE :
					(inData == 8'h0D) ? 8'hD7 :
					(inData == 8'h0E) ? 8'hAB :
					(inData == 8'h0F) ? 8'h76 :
					(inData == 8'h10) ? 8'hCA :
					(inData == 8'h11) ? 8'h82 :
					(inData == 8'h12) ? 8'hC9 :
					(inData == 8'h13) ? 8'h7D :
					(inData == 8'h14) ? 8'hFA :
					(inData == 8'h15) ? 8'h59 :
					(inData == 8'h16) ? 8'h47 :
					(inData == 8'h17) ? 8'hF0 :
					(inData == 8'h18) ? 8'hAD :
					(inData == 8'h19) ? 8'hD4 :
					(inData == 8'h1A) ? 8'hA2 :
					(inData == 8'h1B) ? 8'hAF :
					(inData == 8'h1C) ? 8'h9C :
					(inData == 8'h1D) ? 8'hA4 :
					(inData == 8'h1E) ? 8'h72 :
					(inData == 8'h1F) ? 8'hC0 :
					(inData == 8'h20) ? 8'hB7 :
					(inData == 8'h21) ? 8'hFD :
					(inData == 8'h22) ? 8'h93 :
					(inData == 8'h23) ? 8'h26 :
					(inData == 8'h24) ? 8'h36 :
					(inData == 8'h25) ? 8'h3F :
					(inData == 8'h26) ? 8'hF7 :
					(inData == 8'h27) ? 8'hCC :
					(inData == 8'h28) ? 8'h34 :
					(inData == 8'h29) ? 8'hA5 :
					(inData == 8'h2A) ? 8'hE5 :
					(inData == 8'h2B) ? 8'hF1 :
					(inData == 8'h2C) ? 8'h71 :
					(inData == 8'h2D) ? 8'hD8 :
					(inData == 8'h2E) ? 8'h31 :
					(inData == 8'h2F) ? 8'h15 :
					(inData == 8'h30) ? 8'h04 :
					(inData == 8'h31) ? 8'hC7 :
					(inData == 8'h32) ? 8'h23 :
					(inData == 8'h33) ? 8'hC3 :
					(inData == 8'h34) ? 8'h18 :
					(inData == 8'h35) ? 8'h96 :
					(inData == 8'h36) ? 8'h05 :
					(inData == 8'h37) ? 8'h9A :
					(inData == 8'h38) ? 8'h07 :
					(inData == 8'h39) ? 8'h12 :
					(inData == 8'h3A) ? 8'h80 :
					(inData == 8'h3B) ? 8'hE2 :
					(inData == 8'h3C) ? 8'hEB :
					(inData == 8'h3D) ? 8'h27 :
					(inData == 8'h3E) ? 8'hB2 :
					(inData == 8'h3F) ? 8'h75 :
					(inData == 8'h40) ? 8'h09 :
					(inData == 8'h41) ? 8'h83 :
					(inData == 8'h42) ? 8'h2C :
					(inData == 8'h43) ? 8'h1A :
					(inData == 8'h44) ? 8'h1B :
					(inData == 8'h45) ? 8'h6E :
					(inData == 8'h46) ? 8'h5A :
					(inData == 8'h47) ? 8'hA0 :
					(inData == 8'h48) ? 8'h52 :
					(inData == 8'h49) ? 8'h3B :
					(inData == 8'h4A) ? 8'hD6 :
					(inData == 8'h4B) ? 8'hB3 :
					(inData == 8'h4C) ? 8'h29 :
					(inData == 8'h4D) ? 8'hE3 :
					(inData == 8'h4E) ? 8'h2F :
					(inData == 8'h4F) ? 8'h84 :
					(inData == 8'h50) ? 8'h53 :
					(inData == 8'h51) ? 8'hD1 :
					(inData == 8'h52) ? 8'h00 :
					(inData == 8'h53) ? 8'hED :
					(inData == 8'h54) ? 8'h20 :
					(inData == 8'h55) ? 8'hFC :
					(inData == 8'h56) ? 8'hB1 :
					(inData == 8'h57) ? 8'h5B :
					(inData == 8'h58) ? 8'h6A :
					(inData == 8'h59) ? 8'hCB :
					(inData == 8'h5A) ? 8'hBE :
					(inData == 8'h5B) ? 8'h39 :
					(inData == 8'h5C) ? 8'h4A :
					(inData == 8'h5D) ? 8'h4C :
					(inData == 8'h5E) ? 8'h58 :
					(inData == 8'h5F) ? 8'hCF :
					(inData == 8'h60) ? 8'hD0 :
					(inData == 8'h61) ? 8'hEF :
					(inData == 8'h62) ? 8'hAA :
					(inData == 8'h63) ? 8'hFB :
					(inData == 8'h64) ? 8'h43 :
					(inData == 8'h65) ? 8'h4D :
					(inData == 8'h66) ? 8'h33 :
					(inData == 8'h67) ? 8'h85 :
					(inData == 8'h68) ? 8'h45 :
					(inData == 8'h69) ? 8'hF9 :
					(inData == 8'h6A) ? 8'h02 :
					(inData == 8'h6B) ? 8'h7F :
					(inData == 8'h6C) ? 8'h50 :
					(inData == 8'h6D) ? 8'h3C :
					(inData == 8'h6E) ? 8'h9F :
					(inData == 8'h6F) ? 8'hA8 :
					(inData == 8'h70) ? 8'h51 :
					(inData == 8'h71) ? 8'hA3 :
					(inData == 8'h72) ? 8'h40 :
					(inData == 8'h73) ? 8'h8F :
					(inData == 8'h74) ? 8'h92 :
					(inData == 8'h75) ? 8'h9D :
					(inData == 8'h76) ? 8'h38 :
					(inData == 8'h77) ? 8'hF5 :
					(inData == 8'h78) ? 8'hBC :
					(inData == 8'h79) ? 8'hB6 :
					(inData == 8'h7A) ? 8'hDA :
					(inData == 8'h7B) ? 8'h21 :
					(inData == 8'h7C) ? 8'h10 :
					(inData == 8'h7D) ? 8'hFF :
					(inData == 8'h7E) ? 8'hF3 :
					(inData == 8'h7F) ? 8'hD2 :
					(inData == 8'h80) ? 8'hCD :
					(inData == 8'h81) ? 8'h0C :
					(inData == 8'h82) ? 8'h13 :
					(inData == 8'h83) ? 8'hEC :
					(inData == 8'h84) ? 8'h5F :
					(inData == 8'h85) ? 8'h97 :
					(inData == 8'h86) ? 8'h44 :
					(inData == 8'h87) ? 8'h17 :
					(inData == 8'h88) ? 8'hC4 :
					(inData == 8'h89) ? 8'hA7 :
					(inData == 8'h8A) ? 8'h7E :
					(inData == 8'h8B) ? 8'h3D :
					(inData == 8'h8C) ? 8'h64 :
					(inData == 8'h8D) ? 8'h5D :
					(inData == 8'h8E) ? 8'h19 :
					(inData == 8'h8F) ? 8'h73 :
					(inData == 8'h90) ? 8'h60 :
					(inData == 8'h91) ? 8'h81 :
					(inData == 8'h92) ? 8'h4F :
					(inData == 8'h93) ? 8'hDC :
					(inData == 8'h94) ? 8'h22 :
					(inData == 8'h95) ? 8'h2A :
					(inData == 8'h96) ? 8'h90 :
					(inData == 8'h97) ? 8'h88 :
					(inData == 8'h98) ? 8'h46 :
					(inData == 8'h99) ? 8'hEE :
					(inData == 8'h9A) ? 8'hB8 :
					(inData == 8'h9B) ? 8'h14 :
					(inData == 8'h9C) ? 8'hDE :
					(inData == 8'h9D) ? 8'h5E :
					(inData == 8'h9E) ? 8'h0B :
					(inData == 8'h9F) ? 8'hDB :
					(inData == 8'hA0) ? 8'hE0 :
					(inData == 8'hA1) ? 8'h32 :
					(inData == 8'hA2) ? 8'h3A :
					(inData == 8'hA3) ? 8'h0A :
					(inData == 8'hA4) ? 8'h49 :
					(inData == 8'hA5) ? 8'h06 :
					(inData == 8'hA6) ? 8'h24 :
					(inData == 8'hA7) ? 8'h5C :
					(inData == 8'hA8) ? 8'hC2 :
					(inData == 8'hA9) ? 8'hD3 :
					(inData == 8'hAA) ? 8'hAC :
					(inData == 8'hAB) ? 8'h62 :
					(inData == 8'hAC) ? 8'h91 :
					(inData == 8'hAD) ? 8'h95 :
					(inData == 8'hAE) ? 8'hE4 :
					(inData == 8'hAF) ? 8'h79 :
					(inData == 8'hB0) ? 8'hE7 :
					(inData == 8'hB1) ? 8'hC8 :
					(inData == 8'hB2) ? 8'h37 :
					(inData == 8'hB3) ? 8'h6D :
					(inData == 8'hB4) ? 8'h8D :
					(inData == 8'hB5) ? 8'hD5 :
					(inData == 8'hB6) ? 8'h4E :
					(inData == 8'hB7) ? 8'hA9 :
					(inData == 8'hB8) ? 8'h6C :
					(inData == 8'hB9) ? 8'h56 :
					(inData == 8'hBA) ? 8'hF4 :
					(inData == 8'hBB) ? 8'hEA :
					(inData == 8'hBC) ? 8'h65 :
					(inData == 8'hBD) ? 8'h7A :
					(inData == 8'hBE) ? 8'hAE :
					(inData == 8'hBF) ? 8'h08 :
					(inData == 8'hC0) ? 8'hBA :
					(inData == 8'hC1) ? 8'h78 :
					(inData == 8'hC2) ? 8'h25 :
					(inData == 8'hC3) ? 8'h2E :
					(inData == 8'hC4) ? 8'h1C :
					(inData == 8'hC5) ? 8'hA6 :
					(inData == 8'hC6) ? 8'hB4 :
					(inData == 8'hC7) ? 8'hC6 :
					(inData == 8'hC8) ? 8'hE8 :
					(inData == 8'hC9) ? 8'hDD :
					(inData == 8'hCA) ? 8'h74 :
					(inData == 8'hCB) ? 8'h1F :
					(inData == 8'hCC) ? 8'h4B :
					(inData == 8'hCD) ? 8'hBD :
					(inData == 8'hCE) ? 8'h8B :
					(inData == 8'hCF) ? 8'h8A :
					(inData == 8'hD0) ? 8'h70 :
					(inData == 8'hD1) ? 8'h3E :
					(inData == 8'hD2) ? 8'hB5 :
					(inData == 8'hD3) ? 8'h66 :
					(inData == 8'hD4) ? 8'h48 :
					(inData == 8'hD5) ? 8'h03 :
					(inData == 8'hD6) ? 8'hF6 :
					(inData == 8'hD7) ? 8'h0E :
					(inData == 8'hD8) ? 8'h61 :
					(inData == 8'hD9) ? 8'h35 :
					(inData == 8'hDA) ? 8'h57 :
					(inData == 8'hDB) ? 8'hB9 :
					(inData == 8'hDC) ? 8'h86 :
					(inData == 8'hDD) ? 8'hC1 :
					(inData == 8'hDE) ? 8'h1D :
					(inData == 8'hDF) ? 8'h9E :
					(inData == 8'hE0) ? 8'hE1 :
					(inData == 8'hE1) ? 8'hF8 :
					(inData == 8'hE2) ? 8'h98 :
					(inData == 8'hE3) ? 8'h11 :
					(inData == 8'hE4) ? 8'h69 :
					(inData == 8'hE5) ? 8'hD9 :
					(inData == 8'hE6) ? 8'h8E :
					(inData == 8'hE7) ? 8'h94 :
					(inData == 8'hE8) ? 8'h9B :
					(inData == 8'hE9) ? 8'h1E :
					(inData == 8'hEA) ? 8'h87 :
					(inData == 8'hEB) ? 8'hE9 :
					(inData == 8'hEC) ? 8'hCE :
					(inData == 8'hED) ? 8'h55 :
					(inData == 8'hEE) ? 8'h28 :
					(inData == 8'hEF) ? 8'hDF :
					(inData == 8'hF0) ? 8'h8C :
					(inData == 8'hF1) ? 8'hA1 :
					(inData == 8'hF2) ? 8'h89 :
					(inData == 8'hF3) ? 8'h0D :
					(inData == 8'hF4) ? 8'hBF :
					(inData == 8'hF5) ? 8'hE6 :
					(inData == 8'hF6) ? 8'h42 :
					(inData == 8'hF7) ? 8'h68 :
					(inData == 8'hF8) ? 8'h41 :
					(inData == 8'hF9) ? 8'h99 :
					(inData == 8'hFA) ? 8'h2D :
					(inData == 8'hFB) ? 8'h0F :
					(inData == 8'hFC) ? 8'hB0 :
					(inData == 8'hFD) ? 8'h54 :
					(inData == 8'hFE) ? 8'hBB : 8'h16;

endmodule