module AesMult01Fun (
	input	wire	[7:0]	inData,	
    output	wire	[7:0]	outData 
);

assign outData = inData;

endmodule