module AesBlockMultAlphaFun (
input	wire [127:0]	inBlockNr,
input	wire [127:0]    inTValue,
input	wire [127:0]    outData
);

//TODO

endmodule