module AesMultAlpha02FUn